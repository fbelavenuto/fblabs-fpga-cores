--

LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity teste1 is
	port (
		clock : in std_logic
	);
end entity;

architecture teste of teste1 is

begin

end architecture;
